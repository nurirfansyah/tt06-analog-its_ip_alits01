magic
tech sky130A
timestamp 1713522478
<< metal1 >>
rect 0 630 35 675
rect 15 390 80 400
rect 15 360 25 390
rect 70 360 80 390
rect 15 350 80 360
rect 600 390 665 400
rect 600 360 610 390
rect 655 360 665 390
rect 600 350 665 360
rect 1185 390 1250 400
rect 1185 360 1195 390
rect 1240 360 1250 390
rect 1185 350 1250 360
rect 1770 390 1835 400
rect 1770 360 1780 390
rect 1825 360 1835 390
rect 1770 350 1835 360
rect 2355 390 2420 400
rect 2355 360 2365 390
rect 2410 360 2420 390
rect 2355 350 2420 360
rect 20 315 75 350
rect -55 295 0 305
rect -55 260 -45 295
rect -10 260 35 295
rect 555 260 615 295
rect 1140 260 1265 295
rect 1725 260 1785 295
rect 2310 260 2370 295
rect 2835 290 2895 305
rect 2835 260 2845 290
rect 2885 260 2895 290
rect -55 250 0 260
rect 2835 245 2895 260
rect 15 190 80 200
rect 15 160 25 190
rect 70 160 80 190
rect 15 150 80 160
rect 600 190 665 200
rect 600 160 610 190
rect 655 160 665 190
rect 600 150 665 160
rect 1185 190 1250 200
rect 1185 160 1195 190
rect 1240 160 1250 190
rect 1185 150 1250 160
rect 1770 190 1835 200
rect 1770 160 1780 190
rect 1825 160 1835 190
rect 1770 150 1835 160
rect 2355 190 2420 200
rect 2355 160 2365 190
rect 2410 160 2420 190
rect 2355 150 2420 160
rect 0 0 50 45
<< via1 >>
rect 25 360 70 390
rect 610 360 655 390
rect 1195 360 1240 390
rect 1780 360 1825 390
rect 2365 360 2410 390
rect -45 260 -10 295
rect 2845 260 2885 290
rect 25 160 70 190
rect 610 160 655 190
rect 1195 160 1240 190
rect 1780 160 1825 190
rect 2365 160 2410 190
<< metal2 >>
rect 15 390 80 400
rect 600 390 665 400
rect 1185 390 1250 400
rect 1770 390 1835 400
rect 2355 390 2420 400
rect 15 360 25 390
rect 70 360 610 390
rect 655 360 1195 390
rect 1240 360 1780 390
rect 1825 360 2365 390
rect 2410 360 2860 390
rect 15 355 2860 360
rect 15 350 80 355
rect 600 350 665 355
rect 1185 350 1250 355
rect 1770 350 1835 355
rect 2355 350 2420 355
rect -55 295 0 305
rect 2835 295 2910 305
rect -55 260 -45 295
rect -10 290 2910 295
rect -10 260 2845 290
rect 2885 260 2910 290
rect -55 250 0 260
rect 2835 245 2910 260
rect 15 190 80 200
rect 15 160 25 190
rect 70 185 80 190
rect 600 190 665 200
rect 600 185 610 190
rect 70 160 610 185
rect 655 185 665 190
rect 1185 190 1250 200
rect 1185 185 1195 190
rect 655 160 1195 185
rect 1240 185 1250 190
rect 1770 190 1835 200
rect 1770 185 1780 190
rect 1240 160 1780 185
rect 1825 185 1835 190
rect 2355 190 2420 200
rect 2355 185 2365 190
rect 1825 160 2365 185
rect 2410 160 2420 190
rect 15 150 2420 160
use delaycell_vcro  delaycell_vcro_0
timestamp 1713516147
transform 1 0 5 0 1 -5
box -5 5 580 680
use delaycell_vcro  delaycell_vcro_1
timestamp 1713516147
transform 1 0 590 0 1 -5
box -5 5 580 680
use delaycell_vcro  delaycell_vcro_2
timestamp 1713516147
transform 1 0 1175 0 1 -5
box -5 5 580 680
use delaycell_vcro  delaycell_vcro_3
timestamp 1713516147
transform 1 0 1760 0 1 -5
box -5 5 580 680
use delaycell_vcro  delaycell_vcro_4
timestamp 1713516147
transform 1 0 2345 0 1 -5
box -5 5 580 680
<< labels >>
flabel metal1 0 670 30 675 0 FreeSans 800 0 0 0 vdd
port 1 nsew
flabel metal2 2900 245 2910 305 0 FreeSans 800 0 0 0 out
port 0 nsew
flabel metal2 15 350 20 400 0 FreeSans 800 0 0 0 vcon_p
port 2 nsew
flabel metal2 15 150 20 200 0 FreeSans 800 0 0 0 vcon_n
port 3 nsew
flabel metal1 0 0 35 5 0 FreeSans 800 0 0 0 gnd
port 4 nsew
<< end >>
