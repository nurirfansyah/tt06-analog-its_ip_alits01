magic
tech sky130A
timestamp 1713495731
<< nwell >>
rect -100 260 165 525
<< nmos >>
rect 25 -15 75 85
<< pmos >>
rect 25 280 75 480
<< ndiff >>
rect -10 75 25 85
rect -10 -5 -5 75
rect 15 -5 25 75
rect -10 -15 25 -5
rect 75 75 110 85
rect 75 -5 85 75
rect 105 -5 110 75
rect 75 -15 110 -5
<< pdiff >>
rect -10 470 25 480
rect -10 290 -5 470
rect 15 290 25 470
rect -10 280 25 290
rect 75 470 110 480
rect 75 290 85 470
rect 105 290 110 470
rect 75 280 110 290
<< ndiffc >>
rect -5 -5 15 75
rect 85 -5 105 75
<< pdiffc >>
rect -5 290 15 470
rect 85 290 105 470
<< psubdiff >>
rect -70 75 -10 85
rect -70 -5 -50 75
rect -30 -5 -10 75
rect -70 -15 -10 -5
<< nsubdiff >>
rect -70 470 -10 480
rect -70 290 -50 470
rect -30 290 -10 470
rect -70 280 -10 290
<< psubdiffcont >>
rect -50 -5 -30 75
<< nsubdiffcont >>
rect -50 290 -30 470
<< poly >>
rect 25 480 75 495
rect 25 255 75 280
rect -70 250 75 255
rect -70 230 -60 250
rect -35 230 75 250
rect -70 225 75 230
rect -70 135 75 140
rect -70 115 -60 135
rect -35 115 75 135
rect -70 110 75 115
rect 25 85 75 110
rect 25 -30 75 -15
<< polycont >>
rect -60 230 -35 250
rect -60 115 -35 135
<< locali >>
rect -100 570 165 575
rect -100 545 -90 570
rect -65 545 -40 570
rect -15 545 10 570
rect 35 545 60 570
rect 85 545 110 570
rect 135 545 165 570
rect -100 540 165 545
rect -50 470 -30 540
rect -50 280 -30 290
rect -5 470 15 480
rect -80 255 -25 260
rect -80 225 -70 255
rect -40 250 -25 255
rect -35 230 -25 250
rect -40 225 -25 230
rect -80 220 -25 225
rect -5 200 15 290
rect -70 195 15 200
rect -70 170 -60 195
rect -15 170 15 195
rect -70 165 15 170
rect -80 140 -25 145
rect -80 110 -70 140
rect -40 135 -25 140
rect -35 115 -25 135
rect -40 110 -25 115
rect -80 105 -25 110
rect -50 75 -30 85
rect -50 -55 -30 -5
rect -5 75 15 165
rect -5 -15 15 -5
rect 85 470 105 480
rect 85 200 105 290
rect 85 195 165 200
rect 85 170 110 195
rect 155 170 165 195
rect 85 165 165 170
rect 85 75 105 165
rect 85 -15 105 -5
rect -100 -60 165 -55
rect -100 -85 -90 -60
rect -65 -85 -40 -60
rect -15 -85 10 -60
rect 35 -85 60 -60
rect 85 -85 110 -60
rect 135 -85 165 -60
rect -100 -90 165 -85
<< viali >>
rect -90 545 -65 570
rect -40 545 -15 570
rect 10 545 35 570
rect 60 545 85 570
rect 110 545 135 570
rect -70 250 -40 255
rect -70 230 -60 250
rect -60 230 -40 250
rect -70 225 -40 230
rect -60 170 -15 195
rect -70 135 -40 140
rect -70 115 -60 135
rect -60 115 -40 135
rect -70 110 -40 115
rect 110 170 155 195
rect -90 -85 -65 -60
rect -40 -85 -15 -60
rect 10 -85 35 -60
rect 60 -85 85 -60
rect 110 -85 135 -60
<< metal1 >>
rect -100 570 165 580
rect -100 545 -90 570
rect -65 545 -40 570
rect -15 545 10 570
rect 35 545 60 570
rect 85 545 110 570
rect 135 545 165 570
rect -100 535 165 545
rect -80 255 -25 260
rect -80 225 -70 255
rect -40 225 -25 255
rect -80 220 -25 225
rect -70 195 -5 200
rect -70 170 -60 195
rect -15 170 -5 195
rect -70 165 -5 170
rect 100 195 165 200
rect 100 170 110 195
rect 155 170 165 195
rect 100 165 165 170
rect -80 140 -25 145
rect -80 110 -70 140
rect -40 110 -25 140
rect -80 105 -25 110
rect -100 -60 165 -50
rect -100 -85 -90 -60
rect -65 -85 -40 -60
rect -15 -85 10 -60
rect 35 -85 60 -60
rect 85 -85 110 -60
rect 135 -85 165 -60
rect -100 -95 165 -85
<< labels >>
flabel metal1 -100 575 -75 580 0 FreeSans 400 0 0 0 vdd
port 0 nsew
flabel metal1 -80 255 -55 260 0 FreeSans 400 0 0 0 vcon_p
port 1 nsew
flabel metal1 140 195 165 200 0 FreeSans 400 0 0 0 out
port 2 nsew
flabel metal1 -70 165 -45 170 0 FreeSans 400 0 0 0 in
port 3 nsew
flabel metal1 -80 105 -55 110 0 FreeSans 400 0 0 0 vcon_n
port 4 nsew
flabel metal1 -100 -95 -75 -90 0 FreeSans 400 0 0 0 gnd
port 5 nsew
<< end >>
