magic
tech sky130A
timestamp 1713548907
<< metal1 >>
rect 0 630 40 675
rect 15 390 80 400
rect 15 360 25 390
rect 70 360 80 390
rect 15 350 80 360
rect 600 390 665 400
rect 600 360 610 390
rect 655 360 665 390
rect 600 350 665 360
rect 1185 390 1250 400
rect 1185 360 1195 390
rect 1240 360 1250 390
rect 1185 350 1250 360
rect 1770 390 1835 400
rect 1770 360 1780 390
rect 1825 360 1835 390
rect 1770 350 1835 360
rect 2355 390 2420 400
rect 2355 360 2365 390
rect 2410 360 2420 390
rect 2355 350 2420 360
rect 20 315 75 350
rect -55 295 0 305
rect 470 295 560 310
rect 1050 300 1140 310
rect -55 260 -45 295
rect -10 260 35 295
rect 470 290 615 295
rect 470 260 480 290
rect 550 260 615 290
rect -55 250 0 260
rect 470 240 560 260
rect 1050 250 1070 300
rect 1120 295 1140 300
rect 1640 300 1730 310
rect 1120 260 1265 295
rect 1120 250 1140 260
rect 1050 240 1140 250
rect 1640 250 1660 300
rect 1710 295 1730 300
rect 2220 300 2310 310
rect 1710 260 1785 295
rect 1710 250 1730 260
rect 1640 240 1730 250
rect 2220 250 2240 300
rect 2290 295 2310 300
rect 2290 260 2370 295
rect 2835 290 2895 305
rect 2835 260 2845 290
rect 2885 260 2895 290
rect 2290 250 2310 260
rect 2220 240 2310 250
rect 2835 245 2895 260
rect 15 190 80 200
rect 15 160 25 190
rect 70 160 80 190
rect 15 150 80 160
rect 600 190 665 200
rect 600 160 610 190
rect 655 160 665 190
rect 600 150 665 160
rect 1185 190 1250 200
rect 1185 160 1195 190
rect 1240 160 1250 190
rect 1185 150 1250 160
rect 1770 190 1835 200
rect 1770 160 1780 190
rect 1825 160 1835 190
rect 1770 150 1835 160
rect 2355 190 2420 200
rect 2355 160 2365 190
rect 2410 160 2420 190
rect 2355 150 2420 160
rect 0 0 50 45
<< via1 >>
rect 25 360 70 390
rect 610 360 655 390
rect 1195 360 1240 390
rect 1780 360 1825 390
rect 2365 360 2410 390
rect -45 260 -10 295
rect 480 260 550 290
rect 1070 250 1120 300
rect 1660 250 1710 300
rect 2240 250 2290 300
rect 2845 260 2885 290
rect 25 160 70 190
rect 610 160 655 190
rect 1195 160 1240 190
rect 1780 160 1825 190
rect 2365 160 2410 190
<< metal2 >>
rect 15 390 80 400
rect 600 390 665 400
rect 1185 390 1250 400
rect 1770 390 1835 400
rect 2355 390 2420 400
rect 15 360 25 390
rect 70 360 610 390
rect 655 360 1195 390
rect 1240 360 1780 390
rect 1825 360 2365 390
rect 2410 360 2860 390
rect 15 355 2860 360
rect 15 350 80 355
rect 600 350 665 355
rect 1185 350 1250 355
rect 1770 350 1835 355
rect 2355 350 2420 355
rect -110 300 0 310
rect -110 240 -90 300
rect -20 295 0 300
rect -10 260 0 295
rect -20 240 0 260
rect 470 290 560 310
rect 470 260 480 290
rect 550 260 560 290
rect 470 240 560 260
rect 1050 300 1140 310
rect 1050 250 1070 300
rect 1120 250 1140 300
rect 1050 240 1140 250
rect 1640 300 1730 310
rect 1640 250 1660 300
rect 1710 250 1730 300
rect 1640 240 1730 250
rect 2220 300 2310 310
rect 2220 250 2240 300
rect 2290 250 2310 300
rect 2835 295 2910 305
rect 2830 290 2910 295
rect 2830 260 2845 290
rect 2885 260 2910 290
rect 2220 240 2310 250
rect 2835 245 2910 260
rect -110 230 0 240
rect 15 190 80 200
rect 15 160 25 190
rect 70 185 80 190
rect 600 190 665 200
rect 600 185 610 190
rect 70 160 610 185
rect 655 185 665 190
rect 1185 190 1250 200
rect 1185 185 1195 190
rect 655 160 1195 185
rect 1240 185 1250 190
rect 1770 190 1835 200
rect 1770 185 1780 190
rect 1240 160 1780 185
rect 1825 185 1835 190
rect 2355 190 2420 200
rect 2355 185 2365 190
rect 1825 160 2365 185
rect 2410 160 2420 190
rect 15 150 2420 160
rect 2850 80 2910 245
rect -120 70 2910 80
rect -120 20 -100 70
rect -10 30 2910 70
rect -10 20 10 30
rect -120 10 10 20
<< via2 >>
rect -90 295 -20 300
rect -90 260 -45 295
rect -45 260 -20 295
rect -90 240 -20 260
rect 480 260 550 290
rect 1070 250 1120 300
rect 1660 250 1710 300
rect 2240 250 2290 300
rect -100 20 -10 70
<< metal3 >>
rect 490 310 540 750
rect 1070 310 1120 750
rect 1660 310 1710 760
rect 2240 310 2290 750
rect -110 300 0 310
rect -110 240 -90 300
rect -20 240 0 300
rect 470 290 560 310
rect 470 260 480 290
rect 550 260 560 290
rect 470 240 560 260
rect 1050 300 1140 310
rect 1050 250 1070 300
rect 1120 250 1140 300
rect 1050 240 1140 250
rect 1640 300 1730 310
rect 1640 250 1660 300
rect 1710 250 1730 300
rect 1640 240 1730 250
rect 2220 300 2310 310
rect 2220 250 2240 300
rect 2290 250 2310 300
rect 2220 240 2310 250
rect -110 230 0 240
rect -110 80 -60 230
rect -120 70 10 80
rect -120 20 -100 70
rect -10 20 10 70
rect -120 10 10 20
use delaycell_vcro  delaycell_vcro_0
timestamp 1713516147
transform 1 0 5 0 1 -5
box -5 5 580 680
use delaycell_vcro  delaycell_vcro_1
timestamp 1713516147
transform 1 0 590 0 1 -5
box -5 5 580 680
use delaycell_vcro  delaycell_vcro_2
timestamp 1713516147
transform 1 0 1175 0 1 -5
box -5 5 580 680
use delaycell_vcro  delaycell_vcro_3
timestamp 1713516147
transform 1 0 1760 0 1 -5
box -5 5 580 680
use delaycell_vcro  delaycell_vcro_4
timestamp 1713516147
transform 1 0 2345 0 1 -5
box -5 5 580 680
<< labels >>
flabel space 489 720 540 750 0 FreeSans 800 0 0 0 out1
port 0 nsew
flabel space 1070 720 1121 750 0 FreeSans 800 0 0 0 out2
port 1 nsew
flabel space 1660 730 1711 760 0 FreeSans 800 0 0 0 out3
port 2 nsew
flabel space 2240 720 2291 750 0 FreeSans 800 0 0 0 out4
port 3 nsew
flabel metal2 2895 245 2910 305 0 FreeSans 800 0 0 0 out5
port 4 nsew
flabel metal1 0 630 40 675 0 FreeSans 800 0 0 0 vdd
port 5 nsew
flabel metal2 15 350 20 400 0 FreeSans 800 0 0 0 vcon_p
port 6 nsew
flabel metal2 15 150 20 200 0 FreeSans 800 0 0 0 vcon_n
port 7 nsew
flabel metal1 0 0 50 10 0 FreeSans 800 0 0 0 gnd
port 8 nsew
<< end >>
