magic
tech sky130A
magscale 1 2
timestamp 1713528805
<< metal1 >>
rect 190 6940 29160 6970
rect 190 6860 300 6940
rect 390 6860 530 6940
rect 620 6860 700 6940
rect 790 6860 840 6940
rect 930 6900 29160 6940
rect 930 6860 29570 6900
rect 190 6830 29570 6860
rect 9720 5610 29700 5640
rect 9720 5480 9850 5610
rect 10000 5480 10150 5610
rect 10300 5480 10450 5610
rect 10600 5480 10750 5610
rect 10900 5480 11020 5610
rect 11170 5480 11270 5610
rect 11420 5480 29700 5610
rect 9720 5460 29700 5480
<< via1 >>
rect 300 6860 390 6940
rect 530 6860 620 6940
rect 700 6860 790 6940
rect 840 6860 930 6940
rect 9850 5480 10000 5610
rect 10150 5480 10300 5610
rect 10450 5480 10600 5610
rect 10750 5480 10900 5610
rect 11020 5480 11170 5610
rect 11270 5480 11420 5610
<< metal2 >>
rect 190 7070 510 7110
rect 190 6990 240 7070
rect 330 6990 370 7070
rect 460 6990 510 7070
rect 190 6970 510 6990
rect 190 6940 970 6970
rect 190 6930 300 6940
rect 390 6930 530 6940
rect 190 6850 240 6930
rect 460 6860 530 6930
rect 620 6860 700 6940
rect 790 6860 840 6940
rect 930 6860 970 6940
rect 330 6850 370 6860
rect 460 6850 970 6860
rect 190 6830 970 6850
rect 190 6800 510 6830
rect 190 6720 240 6800
rect 330 6720 370 6800
rect 460 6720 510 6800
rect 190 6700 510 6720
rect 22410 6320 23880 6360
rect 9720 6120 10150 6260
rect 22410 6190 22470 6320
rect 22600 6260 23880 6320
rect 22600 6190 22660 6260
rect 22410 6170 22660 6190
rect 9720 5990 9880 6120
rect 10030 5990 10150 6120
rect 29640 6050 31310 6170
rect 9720 5860 10150 5990
rect 9720 5730 9880 5860
rect 10030 5730 10150 5860
rect 23120 5940 24010 5960
rect 31250 5940 31310 6050
rect 31400 5940 31440 6170
rect 23120 5810 23190 5940
rect 23320 5860 24010 5940
rect 23320 5810 23370 5860
rect 23120 5780 23370 5810
rect 9720 5640 10150 5730
rect 9720 5610 11520 5640
rect 9720 5480 9850 5610
rect 10030 5480 10150 5610
rect 10300 5480 10450 5610
rect 10600 5480 10750 5610
rect 10900 5480 11020 5610
rect 11170 5480 11270 5610
rect 11420 5480 11520 5610
rect 9720 5460 11520 5480
rect 9720 5410 10150 5460
rect 9720 5280 9880 5410
rect 10030 5280 10150 5410
rect 9720 5220 10150 5280
rect 9720 5090 9880 5220
rect 10030 5090 10150 5220
rect 9720 5060 10150 5090
<< via2 >>
rect 240 6990 330 7070
rect 370 6990 460 7070
rect 240 6860 300 6930
rect 300 6860 330 6930
rect 370 6860 390 6930
rect 390 6860 460 6930
rect 240 6850 330 6860
rect 370 6850 460 6860
rect 240 6720 330 6800
rect 370 6720 460 6800
rect 22470 6190 22600 6320
rect 9880 5990 10030 6120
rect 9880 5730 10030 5860
rect 31310 5940 31400 6170
rect 23190 5810 23320 5940
rect 9880 5480 10000 5610
rect 10000 5480 10030 5610
rect 9880 5280 10030 5410
rect 9880 5090 10030 5220
<< metal3 >>
rect 200 7070 500 7140
rect 200 6980 240 7070
rect 330 6980 370 7070
rect 460 6980 500 7070
rect 200 6930 500 6980
rect 200 6840 240 6930
rect 330 6840 370 6930
rect 460 6840 500 6930
rect 200 6800 500 6840
rect 200 6700 240 6800
rect 330 6700 370 6800
rect 460 6700 500 6800
rect 200 6670 500 6700
rect 22450 6320 22620 6340
rect 9780 6190 10120 6270
rect 9780 6060 9870 6190
rect 10020 6120 10120 6190
rect 9780 5990 9880 6060
rect 10030 5990 10120 6120
rect 9780 5960 10120 5990
rect 9780 5830 9870 5960
rect 10020 5860 10120 5960
rect 9780 5730 9880 5830
rect 10030 5730 10120 5860
rect 9780 5600 9870 5730
rect 10020 5610 10120 5730
rect 9780 5480 9880 5600
rect 10030 5480 10120 5610
rect 9780 5460 10120 5480
rect 9780 5330 9870 5460
rect 10020 5410 10120 5460
rect 9780 5280 9880 5330
rect 10030 5280 10120 5410
rect 9780 5220 10120 5280
rect 9780 5090 9870 5220
rect 10030 5090 10120 5220
rect 9780 5030 10120 5090
rect 22450 6190 22470 6320
rect 22600 6190 22620 6320
rect 22450 520 22620 6190
rect 31290 6170 31420 6200
rect 23170 5940 23340 5970
rect 23170 5810 23190 5940
rect 23320 5810 23340 5940
rect 23170 2590 23340 5810
rect 31290 5940 31310 6170
rect 31400 5940 31420 6170
rect 23170 2430 27020 2590
rect 22450 350 22480 520
rect 22590 350 22620 520
rect 22450 310 22620 350
rect 26870 580 27020 2430
rect 31290 620 31420 5940
rect 26870 520 27040 580
rect 26870 340 26900 520
rect 27010 340 27040 520
rect 26870 310 27040 340
rect 31290 540 31460 620
rect 31290 370 31320 540
rect 31430 370 31460 540
rect 31290 330 31460 370
<< via3 >>
rect 240 6990 330 7060
rect 240 6980 330 6990
rect 370 6990 460 7060
rect 370 6980 460 6990
rect 240 6850 330 6920
rect 240 6840 330 6850
rect 370 6850 460 6920
rect 370 6840 460 6850
rect 240 6720 330 6780
rect 240 6700 330 6720
rect 370 6720 460 6780
rect 370 6700 460 6720
rect 9870 6120 10020 6190
rect 9870 6060 9880 6120
rect 9880 6060 10020 6120
rect 9870 5860 10020 5960
rect 9870 5830 9880 5860
rect 9880 5830 10020 5860
rect 9870 5610 10020 5730
rect 9870 5600 9880 5610
rect 9880 5600 10020 5610
rect 9870 5410 10020 5460
rect 9870 5330 9880 5410
rect 9880 5330 10020 5410
rect 9870 5090 9880 5220
rect 9880 5090 10020 5220
rect 22480 350 22590 520
rect 26900 340 27010 520
rect 31320 370 31430 540
<< metal4 >>
rect 798 44700 858 45152
rect 1534 44700 1594 45152
rect 2270 44700 2330 45152
rect 3006 44700 3066 45152
rect 3742 44700 3802 45152
rect 4478 44700 4538 45152
rect 5214 44700 5274 45152
rect 5950 44700 6010 45152
rect 6686 44700 6746 45152
rect 7422 44700 7482 45152
rect 8158 44700 8218 45152
rect 8894 44700 8954 45152
rect 9630 44700 9690 45152
rect 10366 44700 10426 45152
rect 11102 44700 11162 45152
rect 11838 44700 11898 45152
rect 12574 44700 12634 45152
rect 13310 44700 13370 45152
rect 14046 44700 14106 45152
rect 14782 44700 14842 45152
rect 15518 44700 15578 45152
rect 16254 44700 16314 45152
rect 16990 44700 17050 45152
rect 17726 44700 17786 45152
rect 18462 44952 18522 45152
rect 19198 44952 19258 45152
rect 19934 44952 19994 45152
rect 20670 44952 20730 45152
rect 21406 44952 21466 45152
rect 22142 44952 22202 45152
rect 22878 44952 22938 45152
rect 23614 44952 23674 45152
rect 24350 44952 24410 45152
rect 25086 44952 25146 45152
rect 25822 44952 25882 45152
rect 26558 44952 26618 45152
rect 27294 44952 27354 45152
rect 28030 44952 28090 45152
rect 28766 44952 28826 45152
rect 29502 44952 29562 45152
rect 30238 44952 30298 45152
rect 30974 44952 31034 45152
rect 31710 44952 31770 45152
rect 720 44520 17840 44700
rect 9860 44152 10040 44520
rect 200 7060 500 44152
rect 200 6980 240 7060
rect 330 6980 370 7060
rect 460 6980 500 7060
rect 200 6920 500 6980
rect 200 6840 240 6920
rect 330 6840 370 6920
rect 460 6840 500 6920
rect 200 6780 500 6840
rect 200 6700 240 6780
rect 330 6700 370 6780
rect 460 6700 500 6780
rect 200 1000 500 6700
rect 9800 6190 10100 44152
rect 9800 6060 9870 6190
rect 10020 6060 10100 6190
rect 9800 5960 10100 6060
rect 9800 5830 9870 5960
rect 10020 5830 10100 5960
rect 9800 5730 10100 5830
rect 9800 5600 9870 5730
rect 10020 5600 10100 5730
rect 9800 5460 10100 5600
rect 9800 5330 9870 5460
rect 10020 5330 10100 5460
rect 9800 5220 10100 5330
rect 9800 5090 9870 5220
rect 10020 5090 10100 5220
rect 9800 1000 10100 5090
rect 22450 520 22620 550
rect 22450 350 22480 520
rect 22590 350 22620 520
rect 22450 310 22620 350
rect 26870 520 27040 550
rect 26870 340 26900 520
rect 27010 340 27040 520
rect 26870 310 27040 340
rect 31290 540 31460 570
rect 31290 370 31320 540
rect 31430 370 31460 540
rect 31290 330 31460 370
rect 400 0 520 200
rect 4816 0 4936 200
rect 9232 0 9352 200
rect 13648 0 13768 200
rect 18064 0 18184 200
rect 22480 0 22600 310
rect 26896 0 27016 310
rect 31312 0 31432 330
use vcro_5s  vcro_5s_0
timestamp 1713522478
transform 1 0 23848 0 1 5558
box -130 -28 5899 1350
<< labels >>
flabel metal4 s 30974 44952 31034 45152 0 FreeSans 480 90 0 0 clk
port 0 nsew signal input
flabel metal4 s 31710 44952 31770 45152 0 FreeSans 480 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 30238 44952 30298 45152 0 FreeSans 480 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 31312 0 31432 200 0 FreeSans 960 0 0 0 ua[0]
port 3 nsew signal bidirectional
flabel metal4 s 26896 0 27016 200 0 FreeSans 960 0 0 0 ua[1]
port 4 nsew signal bidirectional
flabel metal4 s 22480 0 22600 200 0 FreeSans 960 0 0 0 ua[2]
port 5 nsew signal bidirectional
flabel metal4 s 18064 0 18184 200 0 FreeSans 960 0 0 0 ua[3]
port 6 nsew signal bidirectional
flabel metal4 s 13648 0 13768 200 0 FreeSans 960 0 0 0 ua[4]
port 7 nsew signal bidirectional
flabel metal4 s 9232 0 9352 200 0 FreeSans 960 0 0 0 ua[5]
port 8 nsew signal bidirectional
flabel metal4 s 4816 0 4936 200 0 FreeSans 960 0 0 0 ua[6]
port 9 nsew signal bidirectional
flabel metal4 s 400 0 520 200 0 FreeSans 960 0 0 0 ua[7]
port 10 nsew signal bidirectional
flabel metal4 s 29502 44952 29562 45152 0 FreeSans 480 90 0 0 ui_in[0]
port 11 nsew signal input
flabel metal4 s 28766 44952 28826 45152 0 FreeSans 480 90 0 0 ui_in[1]
port 12 nsew signal input
flabel metal4 s 28030 44952 28090 45152 0 FreeSans 480 90 0 0 ui_in[2]
port 13 nsew signal input
flabel metal4 s 27294 44952 27354 45152 0 FreeSans 480 90 0 0 ui_in[3]
port 14 nsew signal input
flabel metal4 s 26558 44952 26618 45152 0 FreeSans 480 90 0 0 ui_in[4]
port 15 nsew signal input
flabel metal4 s 25822 44952 25882 45152 0 FreeSans 480 90 0 0 ui_in[5]
port 16 nsew signal input
flabel metal4 s 25086 44952 25146 45152 0 FreeSans 480 90 0 0 ui_in[6]
port 17 nsew signal input
flabel metal4 s 24350 44952 24410 45152 0 FreeSans 480 90 0 0 ui_in[7]
port 18 nsew signal input
flabel metal4 s 23614 44952 23674 45152 0 FreeSans 480 90 0 0 uio_in[0]
port 19 nsew signal input
flabel metal4 s 22878 44952 22938 45152 0 FreeSans 480 90 0 0 uio_in[1]
port 20 nsew signal input
flabel metal4 s 22142 44952 22202 45152 0 FreeSans 480 90 0 0 uio_in[2]
port 21 nsew signal input
flabel metal4 s 21406 44952 21466 45152 0 FreeSans 480 90 0 0 uio_in[3]
port 22 nsew signal input
flabel metal4 s 20670 44952 20730 45152 0 FreeSans 480 90 0 0 uio_in[4]
port 23 nsew signal input
flabel metal4 s 19934 44952 19994 45152 0 FreeSans 480 90 0 0 uio_in[5]
port 24 nsew signal input
flabel metal4 s 19198 44952 19258 45152 0 FreeSans 480 90 0 0 uio_in[6]
port 25 nsew signal input
flabel metal4 s 18462 44952 18522 45152 0 FreeSans 480 90 0 0 uio_in[7]
port 26 nsew signal input
flabel metal4 s 5950 44952 6010 45152 0 FreeSans 480 90 0 0 uio_oe[0]
port 27 nsew signal output
flabel metal4 s 5214 44952 5274 45152 0 FreeSans 480 90 0 0 uio_oe[1]
port 28 nsew signal output
flabel metal4 s 4478 44952 4538 45152 0 FreeSans 480 90 0 0 uio_oe[2]
port 29 nsew signal output
flabel metal4 s 3742 44952 3802 45152 0 FreeSans 480 90 0 0 uio_oe[3]
port 30 nsew signal output
flabel metal4 s 3006 44952 3066 45152 0 FreeSans 480 90 0 0 uio_oe[4]
port 31 nsew signal output
flabel metal4 s 2270 44952 2330 45152 0 FreeSans 480 90 0 0 uio_oe[5]
port 32 nsew signal output
flabel metal4 s 1534 44952 1594 45152 0 FreeSans 480 90 0 0 uio_oe[6]
port 33 nsew signal output
flabel metal4 s 798 44952 858 45152 0 FreeSans 480 90 0 0 uio_oe[7]
port 34 nsew signal output
flabel metal4 s 11838 44952 11898 45152 0 FreeSans 480 90 0 0 uio_out[0]
port 35 nsew signal output
flabel metal4 s 11102 44952 11162 45152 0 FreeSans 480 90 0 0 uio_out[1]
port 36 nsew signal output
flabel metal4 s 10366 44952 10426 45152 0 FreeSans 480 90 0 0 uio_out[2]
port 37 nsew signal output
flabel metal4 s 9630 44952 9690 45152 0 FreeSans 480 90 0 0 uio_out[3]
port 38 nsew signal output
flabel metal4 s 8894 44952 8954 45152 0 FreeSans 480 90 0 0 uio_out[4]
port 39 nsew signal output
flabel metal4 s 8158 44952 8218 45152 0 FreeSans 480 90 0 0 uio_out[5]
port 40 nsew signal output
flabel metal4 s 7422 44952 7482 45152 0 FreeSans 480 90 0 0 uio_out[6]
port 41 nsew signal output
flabel metal4 s 6686 44952 6746 45152 0 FreeSans 480 90 0 0 uio_out[7]
port 42 nsew signal output
flabel metal4 s 17726 44952 17786 45152 0 FreeSans 480 90 0 0 uo_out[0]
port 43 nsew signal output
flabel metal4 s 16990 44952 17050 45152 0 FreeSans 480 90 0 0 uo_out[1]
port 44 nsew signal output
flabel metal4 s 16254 44952 16314 45152 0 FreeSans 480 90 0 0 uo_out[2]
port 45 nsew signal output
flabel metal4 s 15518 44952 15578 45152 0 FreeSans 480 90 0 0 uo_out[3]
port 46 nsew signal output
flabel metal4 s 14782 44952 14842 45152 0 FreeSans 480 90 0 0 uo_out[4]
port 47 nsew signal output
flabel metal4 s 14046 44952 14106 45152 0 FreeSans 480 90 0 0 uo_out[5]
port 48 nsew signal output
flabel metal4 s 13310 44952 13370 45152 0 FreeSans 480 90 0 0 uo_out[6]
port 49 nsew signal output
flabel metal4 s 12574 44952 12634 45152 0 FreeSans 480 90 0 0 uo_out[7]
port 50 nsew signal output
flabel metal4 200 1000 500 44152 1 FreeSans 2 0 0 0 VPWR
port 51 nsew power bidirectional
flabel metal4 9800 1000 10100 44152 1 FreeSans 2 0 0 0 VGND
port 52 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 32200 45152
<< end >>
