magic
tech sky130A
timestamp 1713549466
<< metal1 >>
rect 85 20310 10850 20330
rect 85 20165 120 20310
rect 230 20250 10850 20310
rect 230 20165 260 20250
rect 85 20145 260 20165
rect 4890 19625 10850 19640
rect 4890 19470 4915 19625
rect 5035 19570 10850 19625
rect 5035 19470 5060 19570
rect 4890 19455 5060 19470
rect 95 3470 14785 3485
rect 95 3430 150 3470
rect 195 3430 265 3470
rect 310 3430 350 3470
rect 395 3430 420 3470
rect 465 3430 14785 3470
rect 95 3415 14785 3430
rect 4860 2805 14850 2820
rect 4860 2740 4925 2805
rect 5000 2740 5075 2805
rect 5150 2740 5225 2805
rect 5300 2740 5375 2805
rect 5450 2740 5510 2805
rect 5585 2740 5635 2805
rect 5710 2740 14850 2805
rect 4860 2730 14850 2740
<< via1 >>
rect 120 20165 230 20310
rect 4915 19470 5035 19625
rect 150 3430 195 3470
rect 265 3430 310 3470
rect 350 3430 395 3470
rect 420 3430 465 3470
rect 4925 2740 5000 2805
rect 5075 2740 5150 2805
rect 5225 2740 5300 2805
rect 5375 2740 5450 2805
rect 5510 2740 5585 2805
rect 5635 2740 5710 2805
<< metal2 >>
rect 85 20310 260 20330
rect 85 20165 120 20310
rect 230 20165 260 20310
rect 85 20145 260 20165
rect 7510 19995 7570 20000
rect 7510 19955 7995 19995
rect 4890 19625 5060 19640
rect 4890 19470 4915 19625
rect 5035 19470 5060 19625
rect 4890 19455 5060 19470
rect 7510 18780 7570 19955
rect 10775 19895 10835 19905
rect 10775 19855 10785 19895
rect 10825 19855 10835 19895
rect 10775 19845 10835 19855
rect 7680 19750 8000 19790
rect 7680 19240 7740 19750
rect 7680 19230 11700 19240
rect 7680 19170 11580 19230
rect 11655 19170 11700 19230
rect 7680 19160 11700 19170
rect 7510 18770 11300 18780
rect 7510 18710 11215 18770
rect 11290 18710 11300 18770
rect 7510 18700 11300 18710
rect 95 3535 255 3555
rect 95 3495 120 3535
rect 165 3495 185 3535
rect 230 3495 255 3535
rect 95 3485 255 3495
rect 95 3470 485 3485
rect 95 3465 150 3470
rect 195 3465 265 3470
rect 95 3425 120 3465
rect 230 3430 265 3465
rect 310 3430 350 3470
rect 395 3430 420 3470
rect 465 3430 485 3470
rect 165 3425 185 3430
rect 230 3425 485 3430
rect 95 3415 485 3425
rect 95 3400 255 3415
rect 95 3360 120 3400
rect 165 3360 185 3400
rect 230 3360 255 3400
rect 95 3350 255 3360
rect 11205 3160 11940 3180
rect 4860 3060 5075 3130
rect 11205 3095 11235 3160
rect 11300 3130 11940 3160
rect 11300 3095 11330 3130
rect 11205 3085 11330 3095
rect 4860 2995 4940 3060
rect 5015 2995 5075 3060
rect 14690 3025 15655 3085
rect 14690 3015 14830 3025
rect 4860 2930 5075 2995
rect 4860 2865 4940 2930
rect 5015 2865 5075 2930
rect 11560 2970 12005 2980
rect 15625 2970 15655 3025
rect 15700 2970 15720 3085
rect 11560 2905 11595 2970
rect 11660 2930 12005 2970
rect 11660 2905 11685 2930
rect 11560 2890 11685 2905
rect 4860 2820 5075 2865
rect 4860 2805 5760 2820
rect 4860 2740 4925 2805
rect 5015 2740 5075 2805
rect 5150 2740 5225 2805
rect 5300 2740 5375 2805
rect 5450 2740 5510 2805
rect 5585 2740 5635 2805
rect 5710 2740 5760 2805
rect 4860 2730 5760 2740
rect 4860 2705 5075 2730
rect 4860 2640 4940 2705
rect 5015 2640 5075 2705
rect 4860 2610 5075 2640
rect 4860 2545 4940 2610
rect 5015 2545 5075 2610
rect 4860 2530 5075 2545
<< via2 >>
rect 120 20165 230 20310
rect 4915 19470 5035 19625
rect 10785 19855 10825 19895
rect 11580 19170 11655 19230
rect 11215 18710 11290 18770
rect 120 3495 165 3535
rect 185 3495 230 3535
rect 120 3430 150 3465
rect 150 3430 165 3465
rect 185 3430 195 3465
rect 195 3430 230 3465
rect 120 3425 165 3430
rect 185 3425 230 3430
rect 120 3360 165 3400
rect 185 3360 230 3400
rect 11235 3095 11300 3160
rect 4940 2995 5015 3060
rect 4940 2865 5015 2930
rect 15655 2970 15700 3085
rect 11595 2905 11660 2970
rect 4940 2740 5000 2805
rect 5000 2740 5015 2805
rect 4940 2640 5015 2705
rect 4940 2545 5015 2610
<< metal3 >>
rect 8850 22240 10835 22245
rect 8850 22195 8865 22240
rect 8915 22195 10835 22240
rect 8850 22185 10835 22195
rect 8495 22115 10215 22125
rect 8495 22070 8510 22115
rect 8560 22070 10215 22115
rect 8495 22060 10215 22070
rect 8120 21965 9635 21975
rect 8120 21920 8130 21965
rect 8180 21920 9635 21965
rect 8120 21910 9635 21920
rect 7745 21765 9045 21770
rect 7745 21720 7760 21765
rect 7805 21720 9045 21765
rect 7745 21715 9045 21720
rect 7375 21545 8465 21555
rect 7375 21495 7385 21545
rect 7430 21495 8465 21545
rect 7375 21485 8465 21495
rect 8415 20340 8465 21485
rect 8995 20345 9045 21715
rect 9585 20355 9635 21910
rect 10165 20345 10215 22060
rect 85 20310 260 20330
rect 85 20165 120 20310
rect 230 20165 260 20310
rect 85 20145 260 20165
rect 10785 19905 10835 22185
rect 10775 19895 10835 19905
rect 10775 19855 10785 19895
rect 10825 19855 10835 19895
rect 10775 19845 10835 19855
rect 10785 19795 10835 19845
rect 4890 19625 5060 19640
rect 4890 19470 4915 19625
rect 5035 19470 5060 19625
rect 4890 19455 5060 19470
rect 11565 19230 11670 19245
rect 11565 19170 11580 19230
rect 11655 19170 11670 19230
rect 11200 18770 11310 18790
rect 11200 18710 11215 18770
rect 11290 18710 11310 18770
rect 100 3535 250 3570
rect 100 3490 120 3535
rect 165 3490 185 3535
rect 230 3490 250 3535
rect 100 3465 250 3490
rect 100 3420 120 3465
rect 165 3420 185 3465
rect 230 3420 250 3465
rect 100 3400 250 3420
rect 100 3350 120 3400
rect 165 3350 185 3400
rect 230 3350 250 3400
rect 100 3335 250 3350
rect 11200 3160 11310 18710
rect 4890 3095 5060 3135
rect 4890 3030 4935 3095
rect 5010 3060 5060 3095
rect 4890 2995 4940 3030
rect 5015 2995 5060 3060
rect 4890 2980 5060 2995
rect 4890 2915 4935 2980
rect 5010 2930 5060 2980
rect 4890 2865 4940 2915
rect 5015 2865 5060 2930
rect 4890 2800 4935 2865
rect 5010 2805 5060 2865
rect 4890 2740 4940 2800
rect 5015 2740 5060 2805
rect 4890 2730 5060 2740
rect 4890 2665 4935 2730
rect 5010 2705 5060 2730
rect 4890 2640 4940 2665
rect 5015 2640 5060 2705
rect 4890 2610 5060 2640
rect 4890 2545 4935 2610
rect 5015 2545 5060 2610
rect 4890 2515 5060 2545
rect 11200 3095 11235 3160
rect 11300 3095 11310 3160
rect 11200 260 11310 3095
rect 11565 2970 11670 19170
rect 11565 2905 11595 2970
rect 11660 2905 11670 2970
rect 11565 1295 11670 2905
rect 15645 3085 15710 3100
rect 15645 2970 15655 3085
rect 15700 2970 15710 3085
rect 11565 1220 13510 1295
rect 11585 1215 13510 1220
rect 11200 175 11240 260
rect 11295 175 11310 260
rect 11200 155 11310 175
rect 13435 290 13510 1215
rect 15645 310 15710 2970
rect 13435 260 13520 290
rect 13435 170 13450 260
rect 13505 170 13520 260
rect 13435 155 13520 170
rect 15645 270 15730 310
rect 15645 185 15660 270
rect 15715 185 15730 270
rect 15645 165 15730 185
<< via3 >>
rect 8865 22195 8915 22240
rect 8510 22070 8560 22115
rect 8130 21920 8180 21965
rect 7760 21720 7805 21765
rect 7385 21495 7430 21545
rect 120 20165 230 20310
rect 4915 19470 5035 19625
rect 120 3495 165 3530
rect 120 3490 165 3495
rect 185 3495 230 3530
rect 185 3490 230 3495
rect 120 3425 165 3460
rect 120 3420 165 3425
rect 185 3425 230 3460
rect 185 3420 230 3425
rect 120 3360 165 3390
rect 120 3350 165 3360
rect 185 3360 230 3390
rect 185 3350 230 3360
rect 4935 3060 5010 3095
rect 4935 3030 4940 3060
rect 4940 3030 5010 3060
rect 4935 2930 5010 2980
rect 4935 2915 4940 2930
rect 4940 2915 5010 2930
rect 4935 2805 5010 2865
rect 4935 2800 4940 2805
rect 4940 2800 5010 2805
rect 4935 2705 5010 2730
rect 4935 2665 4940 2705
rect 4940 2665 5010 2705
rect 4935 2545 4940 2610
rect 4940 2545 5010 2610
rect 11240 175 11295 260
rect 13450 170 13505 260
rect 15660 185 15715 270
<< metal4 >>
rect 399 22350 429 22576
rect 767 22350 797 22576
rect 1135 22350 1165 22576
rect 1503 22350 1533 22576
rect 1871 22350 1901 22576
rect 2239 22350 2269 22576
rect 2607 22350 2637 22576
rect 2975 22350 3005 22576
rect 3343 22350 3373 22576
rect 3711 22350 3741 22576
rect 4079 22350 4109 22576
rect 4447 22350 4477 22576
rect 4815 22350 4845 22576
rect 5183 22350 5213 22576
rect 5551 22350 5581 22576
rect 5919 22350 5949 22576
rect 6287 22350 6317 22576
rect 6655 22350 6685 22576
rect 7023 22350 7053 22576
rect 7391 22365 7421 22576
rect 7759 22380 7789 22576
rect 360 22260 7053 22350
rect 4930 22076 5020 22260
rect 100 20310 250 22076
rect 100 20165 120 20310
rect 230 20165 250 20310
rect 100 3530 250 20165
rect 100 3490 120 3530
rect 165 3490 185 3530
rect 230 3490 250 3530
rect 100 3460 250 3490
rect 100 3420 120 3460
rect 165 3420 185 3460
rect 230 3420 250 3460
rect 100 3390 250 3420
rect 100 3350 120 3390
rect 165 3350 185 3390
rect 230 3350 250 3390
rect 100 500 250 3350
rect 4900 19625 5050 22076
rect 7375 21545 7440 22365
rect 7750 21780 7800 22380
rect 8127 22365 8157 22576
rect 8495 22365 8525 22576
rect 8863 22370 8893 22576
rect 9231 22476 9261 22576
rect 9599 22476 9629 22576
rect 9967 22476 9997 22576
rect 10335 22476 10365 22576
rect 10703 22476 10733 22576
rect 11071 22476 11101 22576
rect 11439 22476 11469 22576
rect 11807 22476 11837 22576
rect 12175 22476 12205 22576
rect 12543 22476 12573 22576
rect 12911 22476 12941 22576
rect 13279 22476 13309 22576
rect 13647 22476 13677 22576
rect 14015 22476 14045 22576
rect 14383 22476 14413 22576
rect 14751 22476 14781 22576
rect 15119 22476 15149 22576
rect 15487 22476 15517 22576
rect 15855 22476 15885 22576
rect 8120 21965 8190 22365
rect 8495 22115 8575 22365
rect 8850 22240 8930 22370
rect 8850 22195 8865 22240
rect 8915 22195 8930 22240
rect 8850 22185 8930 22195
rect 8495 22070 8510 22115
rect 8560 22070 8575 22115
rect 8495 22060 8575 22070
rect 8120 21920 8130 21965
rect 8180 21920 8190 21965
rect 8120 21910 8190 21920
rect 7750 21765 7815 21780
rect 7750 21720 7760 21765
rect 7805 21720 7815 21765
rect 7750 21715 7815 21720
rect 7375 21495 7385 21545
rect 7430 21495 7440 21545
rect 7375 21480 7440 21495
rect 4900 19470 4915 19625
rect 5035 19470 5050 19625
rect 4900 3095 5050 19470
rect 4900 3030 4935 3095
rect 5010 3030 5050 3095
rect 4900 2980 5050 3030
rect 4900 2915 4935 2980
rect 5010 2915 5050 2980
rect 4900 2865 5050 2915
rect 4900 2800 4935 2865
rect 5010 2800 5050 2865
rect 4900 2730 5050 2800
rect 4900 2665 4935 2730
rect 5010 2665 5050 2730
rect 4900 2610 5050 2665
rect 4900 2545 4935 2610
rect 5010 2545 5050 2610
rect 4900 500 5050 2545
rect 11225 260 11310 275
rect 11225 175 11240 260
rect 11295 175 11310 260
rect 11225 155 11310 175
rect 13435 260 13520 275
rect 13435 170 13450 260
rect 13505 170 13520 260
rect 13435 155 13520 170
rect 15645 270 15730 285
rect 15645 185 15660 270
rect 15715 185 15730 270
rect 15645 165 15730 185
rect 200 0 260 100
rect 2408 0 2468 100
rect 4616 0 4676 100
rect 6824 0 6884 100
rect 9032 0 9092 100
rect 11240 0 11300 155
rect 13448 0 13508 155
rect 15656 0 15716 165
use vcro_5s_taps  vcro_5s_0
timestamp 1713548907
transform 1 0 7925 0 1 19600
box -120 0 2925 760
use vcro_5s  vcro_5s_1
timestamp 1713522478
transform 1 0 11859 0 1 2779
box -55 0 2925 675
<< labels >>
flabel metal4 s 15487 22476 15517 22576 0 FreeSans 240 90 0 0 clk
port 0 nsew signal input
flabel metal4 s 15855 22476 15885 22576 0 FreeSans 240 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 15119 22476 15149 22576 0 FreeSans 240 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 15656 0 15716 100 0 FreeSans 480 0 0 0 ua[0]
port 3 nsew signal bidirectional
flabel metal4 s 13448 0 13508 100 0 FreeSans 480 0 0 0 ua[1]
port 4 nsew signal bidirectional
flabel metal4 s 11240 0 11300 100 0 FreeSans 480 0 0 0 ua[2]
port 5 nsew signal bidirectional
flabel metal4 s 9032 0 9092 100 0 FreeSans 480 0 0 0 ua[3]
port 6 nsew signal bidirectional
flabel metal4 s 6824 0 6884 100 0 FreeSans 480 0 0 0 ua[4]
port 7 nsew signal bidirectional
flabel metal4 s 4616 0 4676 100 0 FreeSans 480 0 0 0 ua[5]
port 8 nsew signal bidirectional
flabel metal4 s 2408 0 2468 100 0 FreeSans 480 0 0 0 ua[6]
port 9 nsew signal bidirectional
flabel metal4 s 200 0 260 100 0 FreeSans 480 0 0 0 ua[7]
port 10 nsew signal bidirectional
flabel metal4 s 14751 22476 14781 22576 0 FreeSans 240 90 0 0 ui_in[0]
port 11 nsew signal input
flabel metal4 s 14383 22476 14413 22576 0 FreeSans 240 90 0 0 ui_in[1]
port 12 nsew signal input
flabel metal4 s 14015 22476 14045 22576 0 FreeSans 240 90 0 0 ui_in[2]
port 13 nsew signal input
flabel metal4 s 13647 22476 13677 22576 0 FreeSans 240 90 0 0 ui_in[3]
port 14 nsew signal input
flabel metal4 s 13279 22476 13309 22576 0 FreeSans 240 90 0 0 ui_in[4]
port 15 nsew signal input
flabel metal4 s 12911 22476 12941 22576 0 FreeSans 240 90 0 0 ui_in[5]
port 16 nsew signal input
flabel metal4 s 12543 22476 12573 22576 0 FreeSans 240 90 0 0 ui_in[6]
port 17 nsew signal input
flabel metal4 s 12175 22476 12205 22576 0 FreeSans 240 90 0 0 ui_in[7]
port 18 nsew signal input
flabel metal4 s 11807 22476 11837 22576 0 FreeSans 240 90 0 0 uio_in[0]
port 19 nsew signal input
flabel metal4 s 11439 22476 11469 22576 0 FreeSans 240 90 0 0 uio_in[1]
port 20 nsew signal input
flabel metal4 s 11071 22476 11101 22576 0 FreeSans 240 90 0 0 uio_in[2]
port 21 nsew signal input
flabel metal4 s 10703 22476 10733 22576 0 FreeSans 240 90 0 0 uio_in[3]
port 22 nsew signal input
flabel metal4 s 10335 22476 10365 22576 0 FreeSans 240 90 0 0 uio_in[4]
port 23 nsew signal input
flabel metal4 s 9967 22476 9997 22576 0 FreeSans 240 90 0 0 uio_in[5]
port 24 nsew signal input
flabel metal4 s 9599 22476 9629 22576 0 FreeSans 240 90 0 0 uio_in[6]
port 25 nsew signal input
flabel metal4 s 9231 22476 9261 22576 0 FreeSans 240 90 0 0 uio_in[7]
port 26 nsew signal input
flabel metal4 s 2975 22476 3005 22576 0 FreeSans 240 90 0 0 uio_oe[0]
port 27 nsew signal output
flabel metal4 s 2607 22476 2637 22576 0 FreeSans 240 90 0 0 uio_oe[1]
port 28 nsew signal output
flabel metal4 s 2239 22476 2269 22576 0 FreeSans 240 90 0 0 uio_oe[2]
port 29 nsew signal output
flabel metal4 s 1871 22476 1901 22576 0 FreeSans 240 90 0 0 uio_oe[3]
port 30 nsew signal output
flabel metal4 s 1503 22476 1533 22576 0 FreeSans 240 90 0 0 uio_oe[4]
port 31 nsew signal output
flabel metal4 s 1135 22476 1165 22576 0 FreeSans 240 90 0 0 uio_oe[5]
port 32 nsew signal output
flabel metal4 s 767 22476 797 22576 0 FreeSans 240 90 0 0 uio_oe[6]
port 33 nsew signal output
flabel metal4 s 399 22476 429 22576 0 FreeSans 240 90 0 0 uio_oe[7]
port 34 nsew signal output
flabel metal4 s 5919 22476 5949 22576 0 FreeSans 240 90 0 0 uio_out[0]
port 35 nsew signal output
flabel metal4 s 5551 22476 5581 22576 0 FreeSans 240 90 0 0 uio_out[1]
port 36 nsew signal output
flabel metal4 s 5183 22476 5213 22576 0 FreeSans 240 90 0 0 uio_out[2]
port 37 nsew signal output
flabel metal4 s 4815 22476 4845 22576 0 FreeSans 240 90 0 0 uio_out[3]
port 38 nsew signal output
flabel metal4 s 4447 22476 4477 22576 0 FreeSans 240 90 0 0 uio_out[4]
port 39 nsew signal output
flabel metal4 s 4079 22476 4109 22576 0 FreeSans 240 90 0 0 uio_out[5]
port 40 nsew signal output
flabel metal4 s 3711 22476 3741 22576 0 FreeSans 240 90 0 0 uio_out[6]
port 41 nsew signal output
flabel metal4 s 3343 22476 3373 22576 0 FreeSans 240 90 0 0 uio_out[7]
port 42 nsew signal output
flabel metal4 s 8863 22476 8893 22576 0 FreeSans 240 90 0 0 uo_out[0]
port 43 nsew signal output
flabel metal4 s 8495 22476 8525 22576 0 FreeSans 240 90 0 0 uo_out[1]
port 44 nsew signal output
flabel metal4 s 8127 22476 8157 22576 0 FreeSans 240 90 0 0 uo_out[2]
port 45 nsew signal output
flabel metal4 s 7759 22476 7789 22576 0 FreeSans 240 90 0 0 uo_out[3]
port 46 nsew signal output
flabel metal4 s 7391 22476 7421 22576 0 FreeSans 240 90 0 0 uo_out[4]
port 47 nsew signal output
flabel metal4 s 7023 22476 7053 22576 0 FreeSans 240 90 0 0 uo_out[5]
port 48 nsew signal output
flabel metal4 s 6655 22476 6685 22576 0 FreeSans 240 90 0 0 uo_out[6]
port 49 nsew signal output
flabel metal4 s 6287 22476 6317 22576 0 FreeSans 240 90 0 0 uo_out[7]
port 50 nsew signal output
flabel metal4 100 500 250 22076 1 FreeSans 1 0 0 0 VPWR
port 51 nsew power bidirectional
flabel metal4 4900 500 5050 22076 1 FreeSans 1 0 0 0 VGND
port 52 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 16100 22576
<< end >>
