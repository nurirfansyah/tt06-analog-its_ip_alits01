magic
tech sky130A
timestamp 1713490626
<< nwell >>
rect -100 260 220 525
<< nmos >>
rect 25 -15 75 85
rect 115 -15 165 85
<< pmos >>
rect 25 280 75 480
rect 115 280 165 480
<< ndiff >>
rect -10 75 25 85
rect -10 -5 -5 75
rect 15 -5 25 75
rect -10 -15 25 -5
rect 75 75 115 85
rect 75 -5 85 75
rect 105 -5 115 75
rect 75 -15 115 -5
rect 165 75 200 85
rect 165 -5 175 75
rect 195 -5 200 75
rect 165 -15 200 -5
<< pdiff >>
rect -10 470 25 480
rect -10 290 -5 470
rect 15 290 25 470
rect -10 280 25 290
rect 75 470 115 480
rect 75 290 85 470
rect 105 290 115 470
rect 75 280 115 290
rect 165 470 200 480
rect 165 290 175 470
rect 195 290 200 470
rect 165 280 200 290
<< ndiffc >>
rect -5 -5 15 75
rect 85 -5 105 75
rect 175 -5 195 75
<< pdiffc >>
rect -5 290 15 470
rect 85 290 105 470
rect 175 290 195 470
<< psubdiff >>
rect -70 75 -10 85
rect -70 -5 -50 75
rect -30 -5 -10 75
rect -70 -15 -10 -5
<< nsubdiff >>
rect -70 470 -10 480
rect -70 290 -50 470
rect -30 290 -10 470
rect -70 280 -10 290
<< psubdiffcont >>
rect -50 -5 -30 75
<< nsubdiffcont >>
rect -50 290 -30 470
<< poly >>
rect 25 480 75 495
rect 115 480 165 495
rect 25 265 75 280
rect 115 265 165 280
rect 25 245 165 265
rect 25 120 35 245
rect 55 120 75 245
rect 25 100 165 120
rect 25 85 75 100
rect 115 85 165 100
rect 25 -30 75 -15
rect 115 -30 165 -15
<< polycont >>
rect 35 120 55 245
<< locali >>
rect -100 570 220 575
rect -100 545 -90 570
rect -65 545 -40 570
rect -15 545 10 570
rect 35 545 60 570
rect 85 545 110 570
rect 135 545 160 570
rect 185 545 220 570
rect -100 540 220 545
rect -50 470 -30 540
rect -50 280 -30 290
rect -5 470 15 540
rect -5 280 15 290
rect 85 470 105 480
rect 25 245 65 255
rect 25 200 35 245
rect -50 195 35 200
rect -50 165 -40 195
rect -5 165 35 195
rect -50 160 35 165
rect 25 120 35 160
rect 55 120 65 245
rect 25 110 65 120
rect 85 200 105 290
rect 175 470 195 540
rect 175 280 195 290
rect 85 195 185 200
rect 85 165 140 195
rect 175 165 185 195
rect 85 160 185 165
rect -50 75 -30 85
rect -50 -55 -30 -5
rect -5 75 15 85
rect -5 -55 15 -5
rect 85 75 105 160
rect 85 -15 105 -5
rect 175 75 195 85
rect 175 -55 195 -5
rect -100 -60 220 -55
rect -100 -85 -90 -60
rect -65 -85 -40 -60
rect -15 -85 10 -60
rect 35 -85 60 -60
rect 85 -85 110 -60
rect 135 -85 160 -60
rect 185 -85 220 -60
rect -100 -90 220 -85
<< viali >>
rect -90 545 -65 570
rect -40 545 -15 570
rect 10 545 35 570
rect 60 545 85 570
rect 110 545 135 570
rect 160 545 185 570
rect -40 165 -5 195
rect 140 165 175 195
rect -90 -85 -65 -60
rect -40 -85 -15 -60
rect 10 -85 35 -60
rect 60 -85 85 -60
rect 110 -85 135 -60
rect 160 -85 185 -60
<< metal1 >>
rect -100 570 220 580
rect -100 545 -90 570
rect -65 545 -40 570
rect -15 545 10 570
rect 35 545 60 570
rect 85 545 110 570
rect 135 545 160 570
rect 185 545 220 570
rect -100 535 220 545
rect -65 195 5 210
rect -65 165 -40 195
rect -5 165 5 195
rect -65 150 5 165
rect 130 195 190 210
rect 130 165 140 195
rect 175 165 190 195
rect 130 150 190 165
rect -100 -60 220 -50
rect -100 -85 -90 -60
rect -65 -85 -40 -60
rect -15 -85 10 -60
rect 35 -85 60 -60
rect 85 -85 110 -60
rect 135 -85 160 -60
rect 185 -85 220 -60
rect -100 -95 220 -85
<< labels >>
flabel metal1 -65 150 -55 210 0 FreeSans 400 0 0 0 in
port 1 nsew
flabel metal1 -100 535 -70 540 0 FreeSans 400 0 0 0 vdd
port 2 nsew
flabel metal1 185 150 190 210 0 FreeSans 400 0 0 0 out
port 3 nsew
flabel metal1 -100 -55 -70 -50 0 FreeSans 400 0 0 0 gnd
port 4 nsew
<< end >>
